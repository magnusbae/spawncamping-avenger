library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity GALProg is



end;

architecture behavioral of GALProg is
begin

end behavioral;

