library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Adress  is

end;

architecture behavioral of Adress  is
begin

end behavioral;

